     TCOPS VECTOR HOLD FILE DUMP PROGRAM VERSION 95.01

     DATE OF DUMP: 12/234/17:42:25.000

     THERE ARE 609 RECORDS IN THE FILE

     THE LAST RECORD WRITTEN IS RECORD 506

     *****  NAMELIST INPUT  *****

      &HFIN                                                                          
       SID=0523401,                                                                  
       ELMSTR=506,                                                                   
       ELMEND=506,                                                                   
       FORM='LONG',                                                                  
      &END                                                                           
1           LONG REPORT OF THE TCOPS VECTOR HOLD FILE                      RUN  1


  SATELLITE ID:    523401                 SIC/VIC:   0234/01
  ELEMENT SET NUMBER:    506
                                          YY MM DD HH MM SS.SSS
  EPOCH TIME FOR ELEMENTS:                12 08 20 00 00 00.000
  START TIME OF FITTED DATA:              12 07 13 16 20 00.000
  END TIME OF FITTED DATA:                12 08 21 15 26 56.000
  RMS OF FIT:                               .128703D+01
  VECTOR TYPE:                            FREE FLIGHT(ON-ORBIT)       
  REFERENCE COORDINATE SYSTEM:            J2000
  CENTRAL BODY:                           EARTH    
  SPACECRAFT MASS:                          .50000000000000D+03
  SPACECRAFT CROSS-SECTIONAL AREA:
    DRAG     .60000000000000D-05          SOLRAD(EPSRPA)   .60000000000000D-05
  AREA MODEL USED:                        BOX-AND-WING           
                                          BOX TOP (M**2)      =   .00000000D+00
                                          BOX SIDE (M**2)     =   .00000000D+00
                                          BOX END (M**2)      =   .00000000D+00
                                          PANEL FRONT (M**2)  =   .60000000D+01
                                          PANEL EDGE (M**2)   =   .00000000D+00
                                          PANEL OFFSET (DEG)  =   .00000000D+00
                                          CRIT. ANGLE 1 (DEG) =   .00000000D+00
                                          CRIT. ANGLE 2 (DEG) =   .00000000D+00
                                          FEATHERING          = OFF
  NUMBER OF ORBS TO GENERATE ELEMENT SET:   3095
  CONVERGING/DIVERGING INDICATOR:
    D.C. CONVERGED                                                  
  ORBIT THEORY USED:                      COWELL                 
  ATMOSPHERIC MODEL USED:                 JACCHIA-ROBERTS
  CARTESIAN COORDINATES:
    X        .42164000000000D+05 KM       XDOT       .00000000000000D+00 KM/S
    Y        .00000000000000D+00 KM       YDOT       .30746662829706D+01 KM/S
    Z        .00000000000000D+00 KM       ZDOT       .00000000000000D+00 KM/S
  KEPLERIAN ELEMENTS:
    SMA      .42164000000000D+05 KM       LAN        .00000000000000D+00 DEG
    ECC      .00000000000000D+00          PA         .00000000000000D+00 DEG
    INC      .00000000000000D+00 DEG      MA         .00000000000000D+00 DEG
  SOLAR RADIATION PRESSURE COEFFICIENTS:    MODELING IS ON         
    CSUBR    .14000000000000D+01
  DRAG COEFFICIENTS:                        MODELING IS ON         
    CSUBDZ   .20000000000000D+01          RHO2       .00000000000000D+00
    RHO1     .00000000000000D+00          RHO3       .00000000000000D+00
  THRUST MODEL COEFFICIENTS:                MODELING IS OFF        
      .000000D+00     .000000D+00     .000000D+00     .000000D+00     .000000D+00
  RIGHT ASCENSION:
      .000000D+00     .000000D+00     .000000D+00     .000000D+00     .000000D+00
  DECLINATION:
      .000000D+00     .000000D+00     .000000D+00     .000000D+00     .000000D+00
  JOB ID:   user                          SYSTEM:   GTDS    
  MACHINE TIME:                           ** 08 21 13 26 22.000
  MACHINE ID:                             us
